module global_params();
    parameter DIG_CTRL_V_WIDTH = 12;
    parameter P_GAIN = 100;
    parameter I_GAIN = 5;
     

endmodule